* C:\Users\PREZENS\Desktop\CSE250\LAB 2\Schematic1.sch

* Schematics Version 9.1 - Web Update 1
* Fri Nov 20 22:53:35 2020



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic1.net"
.INC "Schematic1.als"


.probe


.END
