* C:\Users\PREZENS\Desktop\CSE250\Schematic1.sch

* Schematics Version 9.1 - Web Update 1
* Mon Dec 21 15:03:10 2020



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic1.net"
.INC "Schematic1.als"


.probe


.END
